module Float8E4_pack(
    input [31:0] f32_in,
    output [7:0] f8_out
);






endmodule