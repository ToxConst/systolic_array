module Float8_unpack #(parameter E = 4, parameter M = 3, parameter BIAS = (1 << (E-1)) - 1) (
    input logic [7:0] fp8_in,
    output logic [31:0] f32_out
);








endmodule

